`timescale 1ns/1ns

 module System ( reset2,clk, rst, sw_0, uart_rxd, 
 a_to_g, AN, DP,led1, final_output1, reset, hsync, vsync, rgb, sw_1, BTNR, BTND); 
  
  //parameter image_size = 11*11, weight_bit=4, output_bit=4, input_bit=1,hidden_layer=30,out_layer=10;
  //parameter image_size = 11*11, weight_bit=4, output_bit=4, input_bit=1,hidden_layer=200,out_layer=10; //Attempt With 200 Layers
  parameter image_size = 11*11, weight_bit=4, output_bit=4, input_bit=1,hidden_layer=100,out_layer=10; //Attempt With 100 Layers
  input wire reset2;
  input wire BTNR;
  input wire BTND;
  input clk;
  input reset;
  output hsync;
  output vsync;
  output [11:0] rgb;
  //input wire clk3;
  input sw_0;
  input sw_1;
  input  wire rst;
  input   wire        uart_rxd; 
  wire [(image_size*input_bit) - 1:0]input_features0; //define the input features (121 dimensions by 1 bits) 
  wire [(image_size*input_bit) - 1:0]input_features; //define the input features (121 dimensions by 1 bits)
  output wire [6:0]  a_to_g;
  output wire [7:0] AN;
  output DP;
  output  led1;
  //output wire clk3; 
  output reg [output_bit-1:0] final_output1; // to distinguish among 10 different digits
  reg [output_bit-1:0] final_output; // to distinguish among 10 different digits
  parameter WIDTH =   7;
  //topology: 121:30:10
  reg [(image_size*hidden_layer*weight_bit)-1:0] weights_NN1_layer1;
  // initial weights_NN1_layer1 = 14520'hfedde0201111ede0440f021f01022fe021001121def13110132e0d12210fefdfee10042242fdf0ef224441effdd024412f00dde042f0f00eddf10ef0000ee0ff2310fedd1fd120f1fef1fe30df1fef43241df10e33224eeefff0fde4eddfed1fe22fdd1ed122320ed0dd242201fe1ddf22ff1000fff0100100000f0f0321001d0f03332011f1ef4232f0101e03201e200eddddddd22edde2f01d2300e14432d231ee34221d110de211fff0000f2211f0000000ff0000fdddd041110dddddd1231fdef1fd02101100eede0e0f0f000020de220234441ed222202420dd1111ffddddd00000fedddf0effe0feef00dde000f00011000ffedf0121f0eeff0e031def00f1f021de034230dfdd0f2421200004eddd030f420fddef2e2421ddef11f2121dde0100210fddf0000211000000002233310fe00144300fef2e2331feff03d0430ddef23e040dddf102ff400dd01120142fffdf13f24131ede02013330ddf2101323fdd000010000000000011fde2010010ffde120100f0ff01ff102f0f0010ff2111def4f1f12420d04f000240edf3020042fdd021000230dd22200022edd131000110001100000ff0feddf0010f10ff10f02f0000144110f00344442fff1213fd13f000feddde0f0f01fdf0dee0f00ee11fd0100fde21fe12210ef000010211000000ff143334111e032320fdf3f2211f0fd23e132f01fd34f13fe11ed24f23f201dd04f141032dd13d24ff32ed13d14201fff32f13301fef110011000ff000fddfffdef0fdf11101feff001342100f1013433310f00120e133ffeffded1220011fdf12ef1110ed14fdf2110ede2de0202ff011f02201012111221011210edddf02ef00f0ded11ddf021efd11ddf231ded2dde2342d1e1dd1444213d2ddf222110d1edd32311ee11ddf331ede00ede11fde00001110fff000110f0fdee0ff1000fedd0df1021effd0dd1012ff1f0ef1f12112110f3310ee4121f111fdd42310d10dde34222dffdde241221ffddd1200121000f000f00234fef20edd04300f12fdd1431fde2fef241ffdf1dd24414edf0dd23413ddf0dd2f244ddefeef0340ed01eef333ef020fef341de0100000000000000000fdddf01000f0ddd22000014dde4011f0111df421120000df43f00ff0fd41410ff01013200fde10110ffeffef0120df11f0e130dd0000000feef00f00f0131d0ff11f2242feefffdf1440ef0eeeee3430f001ddd144121fdd112e1234fe1ef3e211430ff0fef01341fe00fe002320020ff000ff0f000000fddff02ff0feeefe020e0deddff11ffffeee0f0100ffff1422200e0fff344ef1ff1ed44ff00f24fdf4011ef230ddef20f0221edff0000111000110000ff0000ef00ef0ffefd1100ffef20f0f21fff0fddff200f0111de2311f24430124100343df21300443ddf001f222fde1ff0141ffdd01000122000110000f000ff1000fff01111e000de01ff101fedf23200e11fe143fffe020242dd12e01044fdf42f1000ddf1311110eded011200edeedf0010ffff00f0100113411243000330ef1311f031fe023430f0000e2324310110edf0241200dfdd123130242f22220431011433104400012320e341ff111f00100ff000f001221ff4420032101e341f021021d24000ff231f242010011d00221210edeff2302000e14f12f1e1f011032e1f02322020f0023131000f0000000ff001fffffffff010eee02feef3100df00ff0321ff020e0f2120000102f10333e01210ef44ddff100de0ddf110f0fddddf31000fddde0420f0ffff001100000ffe0fdde0210edf1de01101ee240e1010ff0232010f00ef11e0f1e0fd341e000e014421000fef344121fe0efeff110de0efede13fdf0ffeef00ff0002211ff02402320ef0e130230ff21ef11220f23eef1f101244fde1e0ef344dde0e0ed4310fe1dfdf3131fd2eeef1221ee1fef0f12fd110000000fef0010f1200fff0111111021f012100211ef101124212e1101234310e220112441f1311022442f13011fe21fe020000021ef11ff0120ee001000001000f000fef0fffee001010ff0fd00221ff120f0100000213f021fed0124e040eddff440240fefde34022f0dfde2412101ed0f11002110ef021001012101111011331ddd2100143fddd310f043fedf200ef322fde3f1ee2300d02f0ff0022d20f00e0022d0f00e0122fe0001ff230fe0f00f0221ddfe00011100f0f00000210143101343fde12200441dddf0311441ddde041143dddd0131341d1441143343203fdf33234000ede32133ee0df0210320edd011011110f000001221fdfe0f03200dff14fe3020e1f140d1f00ffd141d0e11e0dd41dfff100dd430fff10fdf22200f01ee013211f11eeff210f121ef0ef00001000ff00010f021ddd10ee0334fee2fe002242ef2fe023231ff20f232e0f002ff12dddf101ff130df21f2fe042d121e21ef441221011ee243110000feef011100feedef234101ffedf03400210ef02441e10eff12441e20e0f32230e30df134331e31dddf4422e40ddde2130e22fdd1211ef10fee23120000001221110;
  // (200 Neuron Attempt) initial weights_NN1_layer1 = 96800'h0001100100001100011100000ff01010011fff0000ff20ff000fddf2010100dde000111110f10f0100133220f00000001000000f00000000000000000000001fff00f00000ef000e0ff00ef0f0efef010111ff0df112111001112edd00f00212edd110f0021dd02200002fdef12010f0fdef010000000f0000011121edef00f0120ef0f00df001000f0ede243200f0edf44220ff0dd010210fefddff0121feffeff03110f00ef0231ff000ff211eff00000000f00000010000110001000000000100000000000f0010000011000010010100000f0f0000f01000001000000000110000000000000000000000000000000000000fff000f000ffe0100f00ffef0101001ff00010200000000ff4f0000010ff2e00f010e000e00f00f011ef010f0f00fef00fffff00f00000000000000000011f000001111100010000111100100011000001011111001010100f0011000100110000001011100001010110000100000100001000000000000000000fff000100000f01001001001331010001221000110110edd00000000dfff00f0110020f0f000fef10f00010edf01001100fff10000000000000000f00f000000f0001110000f011110f00ff110000f0100121001f010011f001f000011ff00000ffeff0110010ffff011101ff0ff010000010000000000f01220ff0ff011211fe0f001fff10f0f21ffff110101fe01f2001110efe02011110ddd01f11112ed04f0110112132ff110011010ff10000000000000000000121001000f01100f000fe0110f0000f01021f110ee002310200ed013210210fee12210110eef01200111eef012000110ef111000000000100000feff01000feddddf1100edddedf22f0edf00e021f0e02310f21e0120123121ef220000f11ff20ffffff0ff10ffefeffe010ffffff0f00ff00000000000000011000000000110f010f00011000000111100f1000101100f10f0001101e1ff0001011e1ff0f00010f10f0000000f0000000010000000000000000010ff00000011ff0100001210f0000002120ef0f0000111ef1f0fff112df1f0fff021d11f0ff002fd1100ff011ee100000121ee0000001110000000feeef022100eeeef01100fffeff0220f0ffff0111fe10e0221000e10e0232110e01ee011110e00fde11120f000dd0011f000fed00010000100011000000000fddf010100deddf01010eedddd01110f003edf001ff0322fff00f0241220e0112100011000220fff110fff00ff01000ffffff110000000000000000000ff00110001100f00010111100100011110001000f011f200000ff00f200100100001001ff0110000010f011100100f011100010000000000000001000110001000ff011000f00001110101100110111000ffeff001110ff0101011000100110010f00ff11000100fef11001100ff0100000000000000110011eef00001122fef10f012210ff1ff1220f0f01ff1110e0f01ff011feff01ff111ff00f1f0113000f0100012110f00f000210100000ff0000000000f00023100ff0000111000f000011000ff0100110010fff10010f10ffff0000f10fff22110f1fffe12110f000ff01010f0000f0101000000000000000011feef0001111fede0101110ffee110111f02ee12f012024fe22f00f1430e12f11ed120f21001fe00ef11001000ef0000011feef0000011000f0000001110fff00011100000000000000f0000000ff000000010f01000f0002201100f1001201001000010110000010000000000100001000000000000000000000fef0000000fffff00000ff00f00010ff010000000f0110100001001e0310000f00de3210f0f1fdf21000011dd01001000fef00000100000000010f000000000001121110001112420100112420ffff01120ddd0fff0efef0010000fff00000010ff00010100ff1110ff100000110000000000000000000000000f000110f000f00000f0000ff100000001ef10ffff023ef1f0f01043f010f00ef220100000ef21000000ff011000000ff111000000000100000000000f00000110000f0f000100000000001000000000000011f0000ffff11f0100ffff110010000ff011110000fe011010000ff01000001000000001110000f00111000000001000001100000011f0000101110ff0000010000ef100000011f0101f010110001100100000010001000f00000001000000000000000000ffff00fff00f00111ff11000000ff111011000022f0011114221ef0001100feef0f000fef0f00000fff01000100ff00100000000000000000000011000ffff111100000ff0111001000000110f10000ff110f10000f020f00000fd120f00000ef11ff00000ff10f00000ff0200000000000000000ff0f01ff00f0ffff1ff0fffff000ff0ffff1101000ffff12100ffff0df44ff0ff20d040000f041dd20100f121ddf11000111fefff000001000000000000ff011000000fef00100010ef10020111ff0000200110010f02101ff230f00110e01100f0010f00100f0001100110ef00110f00fff0000000ff000011000001001100f0100001000011000000f000f00000f010eef0000000f00000000f0110101000121111100011111110f0f0000110ff000ff000000001100fffef00010fe0fff0000fef111ff00fff0003ff000fe0f040f000ff1e041000f000f02000000000f000000ff00ff0000ffff0000000000000000000f0fff1100ffffedf1000fef0ddf1f000ff00de0e0011232e11f01233000410f0fefff10feffed12200ee0fef110feff00f0100ff00000000000000000000ff0100fef10001000fe022110f00fe032210ff100221100ef00000ff00ee0fef0ff1fee0edf10010ff0ed0111000f1ee0110010000000000000001100121000121fef01100221eef0120132fefe0021120efef001123ff1210021221110ff0211110ffff010111ff0f00000210fff00000011000000000ff00012100ffff0001100fffffef000110ff1fffff1000121ff0f000112110fe000100220fe00010111fef000000ffee00ffff00fff00fff000000000000000000100fff00010000ff010f10000000000100010121f020f0ff131f0001fe01100fff1ff11101ff00011121fef00000000ee00000000ff00000011111110f0001100010f0001000f00000010feef00011102ee0000012330f0000012300ff00f0110f001001110ff011001000ff0100000000000000111111fff001122110f00f1121ff0f01f120fefff01f010eefff010020ffdf011f121fef0001f0200000f010011210ff000112210ff000000000000000010001110011000000100100000001000000000f000010000ff100000110f00000001100f0000001100f00f00011000000000000f000000000000000000000fff00000100fef0100110ffde0000110f0ddf00110f010de0f0001332f00fff0f01111f0fffff1111000fff011100fffff11010000000110000000000f0000000f0fe0001000f0ff000100ff0fe011000000ff101ff112101101ff21fff1200f0010f010f0f0000011ff00000f010f00000000000000000001221000000001110f100ff0111f0000ff01110010ffef010011feee0110f110fef11110011ee000000012fe00001001100010000001000000000000000fff0001010000f0000001111f0000100121011000f01f11110ffffff21110f0000021100000000111000f000011010010000100001100100000100000011001100000001000001010010f0110000010f110f0f1010010fff01f0110000101000000011011000001110110001111000000000000000000eef0eef000eef11fff11fff1320fef0f0f22110de0f0010e1feffef10ee2201ff030f44ff100000340def00fef11ddff00fff00f000000000000000001100100001110f01fe01110ff010e0111ff00f000100012fe0f0100123eddf01e02331ef010ff101220010ff001200000ff000110f000000000f00000000100f00000ff000ff0f0000000ff0ff00000ff000011100000100421ef1001ff20eeef001fff0fef01010fffff0121000ff0f001000000000000000110f011000010fe0110f010fff0110f1000f00100f10f0001001f10f1220012000000fef1110110ffef110012ffeff0001110feff000001100000000000010000000000000000000000000010f011ff00010f1100f01f10000f0f01e0010011011f1000010f100100100ff111000000ff10000000000000000000000000ff001001100fff010011000f001001ff010000000ee011210f00ff01011ff00011000fe001111000ffff0110000fff00100000000000000000000000000000010f010010f010f01000f00ff000f01021ff001f01022f00f0ff0111f00f0ff011110ef0f011010fef0f010100ff000000000000001100101100000001111000ff011001000ef110f00000ff121f01000001ff0010010f0000101010f0010011011000f0011000000f0000000000000000000f00000100fff00f0010ffff000010fffeee0100fff0ef211100e0010332100f121ff010110130fe000000110ff0fff00110fff00000000000000000110ff010000100ff1121f0000f01120e000ffff120f0f00fef12000010f0011010f0f11010000f0001100000011010000001111000f00000000000000000110fff00010210f0f00000110fff0ff11000ff01ef200110001ef40000f0f1df40f0ff001e041e0ff001f031e0ff01100221ff001000111000000001101111000011001221ff00fff0211ffff0fff222f0feeff0123120edf0ee021121111ee00112200fef1001220ffe000002200fff0000110000000000010ff1000111feff0000010fef002000010ee2110120feefeddd0321fefff00f23220f2342f0110ff2121f0ffee010100fffed0110f000f00000000000000220f0ffff1f240efff000d04fdf00100f04fdf00001134fdf00001013efffef110feef00011110f110101ff00f1110ff000f01100fff0000000000000ff0100100f0012200100001233110000222021100f11fddf1100f01fdfef100011002ef0100f0f11ff0110fff110f0110000010000000000000000f00011000ff000111000000000110000f0100110010f0001010010ffff0110010fff001100100ff000100100ff001100100000100000000000000000000f00110011ff0000101100f01000010000000fff100120fdf0f1fe132fe00f1ee0110001f1ff0110001f00ff11000000000010f0000000000f000000000ff00011110fedf01111101fe011ff0123fd101ff0122fd001fef001ef100ff010200000fff110000f00f011100ef00f01110ff000000000ff000000110ee00000f00fdd1000ff01eef101ff001234400fff114410000fe1feddd0ff1110ddddff00101110000000000000011ff00ff000000000000000011011010001100010000000000000110000100001100110fff011010ffff0000010110f00100000011111000000011110f01001100000000000000000fff0edef01fffff0f0f01f0fef311f1100ff2400f11000041f0f1001032ef1f10f022fe000100f1fe11ff1000ff011f0000fd00100000111000000000000000000001001000f00011111100000011011101000001111011000f010110001010100000010110110000111100010000101000000000000000001100fee0100221f0ed011020f11fd0200210011e120011fff0f110f12dfe0f11f022dffff210032ddfe0120022fdee1110122fef0110001110001000000000111100000011000000001110001000011000011000120000110000f0001000010f00010000001001100100101011000000010000000000000000000110f000f000100ff00000001ff000101000ff11001010020f0000003410ff000f132e0ff0ff021ef0000f0010ef001001010ef010000000000000000011ff0100f0121eef20000120dee00ff0210e0010ef121f33120ef112f1fe00ef10f10ddf0f010020ddf0f01121fef00000131ef01000111000000000110f0000011110ff0000101211e0000f01121e0010fff032ff0100ff022f000001de110000001fe0101100010fff01000000fff100000000000000000000fddf000000fedee010000effff0001001320ff001012311fff0011100100ff1210ff01100f0f0ff010010efff0010100ffff011001100001100012222feef0012220fedf1f0210fffef1ef310fefe12de31ffeff02ef211feff02ef4221e0f02f12230d0002f1121fd0f0101100eeff00010000000000000000000000000011100010ff010010100ff0111101100111001010f111fff001ff000f0ef010f01000ff0000010fff00001100f00000000000000000000000000000f000f0000000010f000000000ff000001100f0100001120010010010fd010000000fff00000000ff00000100fff0000000000000000000f00f0110000111ef1100f1110ee1100f1110ff110001f0ee010f13ed2100f0f33dd220f01f32dd22ff01f21edf1f001011fe0200100001000000000011010101000000000e010100110fe010000111ee010011111ee11f012310de11ff11111fe10ff000010000ff0111000010f00110ff000000000ff0000fff00fff00f0011110f00f0011210f00f010110ff00f10f11f1f0001000f02f00f000ff10010ff00f0011100f00f011100f001000010000000000000001000000000000f0110ff000000000ffff000010100ff00010110100001fe110100010de11100011fdf00001110eeff0011110eff0000010000000000110001100011000f1100000010001000f01100101000010f00110100fffff11011f00000010000001001100010000011000010000000000000000000000000110000000001000100f000000f10f0000110f1000011110f1000011110f10fff01110f1ffff01110f00ff00110000ff00111000000000000000000000220010fff01120f10ff00011f0100010022ff1ff00f012ef100fff011fe0000012100f0ff0f1220ff00011111fe00ff00110ff00fff000000000ff0f0020010ff000130f1fff00023e010f011033df0fe00ff22ef000fdef11ff00f0f0210ff0ff002111fffff111110f00ef011110f00fff00000000100011110011100f0111011100ff00211110fef00111220ffe0101110ff0ff0111210010ff11111000ff021011000e011001101fe0100011000000000000000110000000100100000001001000f0011101100000000f011100fff0001011f000011101000000010000000010000000001100000000000000000110ff00000110feef10000000f0000f0100f00010f1000f11110f000111021000010fdf11110120edf01010031ddf01000120ddf110001110001000000000001000ff01000000000011001000ff02111000000111100f0000000000ff10ef00000f01fef00001000fef01001100ff00100100000000000000000000000000000110000000011100010f0111100110f0000ff110000ffff011011f00011100100001000001000111000000001110000000000000000001000110001110ff01100221feff1101220efef010120efef001022ff02100112201100f0102110ffff010111ff0ff0000110ffff000000000000000000ff0f0101110fffff012221000ff021121220df011112330e0010f0322ff101fef100f01010ff100ff00100f00000000000000010000011010000000100f01210010ff00000010000000000000010010001000121000000010f100100001001001f00000111110000000100000f0000100000000000000000011111ef00000111fdf10ff0112ed010f01002dd12f00f113ed22f021112ee12e041f0fef22f131dffef11f021efef1110011fff01110011000000000000f011100000000110f00000001100000010111001000000000f0fffff0000f0ff0001000f0ff0000000f00f0010000f000001000000000000000000000110000000002111000fff01210010ffe021ff010f0011ef00100001ee11f110f02ff000011110010ff0000000100000000101000000f0000000000000100f0000ff0110ff00ff02310ff00001321100010133ff00ff0022feeeff0f0fde0ff010ffed01f0110000010ff1100f001000100000000f000000000000f0010100000f010010f010f1100000f00011e010110f000f000120f0f0f0012100ff0f0011110f010000110fe010001110ff000000000000000000002100001010000100001fff0110022fde10110131eeee11002210fdd31001210fd011011200fe22100121fef22200011fef12100000000010000000000f000000ff01ff01100f011ff011100110ff01101121fff01001220ff0f1ff120ff00f1ff0f0110ff1ffff11100010fff00000000000000000000010100000000ff0110000000f00100000000001ff011000000ef001221fffe0101320000f10f0fee011110fffef001110ff0f000000000000000000000f0000000000ff1ff000100001ff000100010ff01100121fff11010231d000000f21de101000f0eef0100000ffff1100000ffe010f00000000000000110000fff0011112100000011111000000122ff00000010eddef01f0f00fe000100120ff0001ff222f00f000f12320fef0f1012100f0000ff000000000f0110121000f110f10102211fe101102200e02100f00000101fef0ff0ed00def00fdde43eff11fde441ff00fee0421f001fef12211000000000000000010ff000001110fe00f000110ff000001110f010100100f020120000dd32f021110de110f11111de000f00111fe000f0001110ffff000011000f00000ffff010100ffffee01100eff0ed01000f001fd12ff0e0fff032eef0100222edd0022130ddde0010f0eeeef0000000fff00000000f0000ff0000000000f01000000f00010f0100f00010011000111100100011000010f0010ff0001f01100ff0100f00f0fff0f0010ff000f0110100100f011000000000000000000f00f011f0fff00f010fedef000011fd032001000f0431000f0f032ef00f00f33ee110ffff1fe021ff0ffef0010f000fffff0ff000000000f00000feefffef000fee01110f1110f133210110011124410001000f2420000ffdde420110f0fdf220100fffe011001ff0e000000000ff0ff0000110000000011000ff000001100ee010011100ed01ff11000de11f011101ff11f0121210f01f011f0ef01100110ffff0100110fef00101110ef00000111000000000000000ff0000000110ff0ffff11210f00ff000131f0000f0fe320100fffef11111ffff0001101000f000011110ff00000000000000000000000000000ffeef00000fdffeef1110ef000de130001100ed21f000001ff20e10e0012310d10021244fed0001ffedddef0010eddde0fe00fffff000eef0000000011000feef01100fffeee0000fefeefe0f0fde20e0f1e0ef3210111ff133000101ef21ffe0001ff011f10f000fdfff000000fefff0fff0000000000000012111111001210f00f110111ef00f110110fff0f11f0110ffff11f100321001111111300f010120000ff11f12000f0010f1210ff00000100000000000000000000000001000f000000001001000110000010011110000101000000000000010000000000000100100000f000000000000100000000000000000000000001110000000000000000000000010000000000f0001000000f00f100000010000000000010000000000100000000101000000000000000000fff0011000ffff011100fffff01110ff0ffe0000ff00ff1100f0e00ff321f00e01fe221010f12fd02111ff110de0010f011fee000000001000000000000100110000000f0110f00f0000110f0ff021121ff1f011f011fe10ffff011fe10f000111fe1fef00000ff1ff0110000f1ff010f00000000000000000000111f000000111fef100000010e010010ff1ee11011f000ff110110100ff11f021000f0110110ff00001f000ff000110000000000000000000000000001100000000011100000ff01101000fff00f01100f0000ff111000000f1ff110ef1001f000112101000000110f00000010000000000000000000000000011110ffef0012000ffe00f01ed0fff020ffddf000f101ed000001421422021223ff222f11230ddf00001210effff0100ffef00f000f000000000fee00111101fe011100011000010ff0121f0010ffff410001001ff1100fdedefeff02132feeffef124430ffffe012321f00fff02200f00fff010f000000fffffef00fff000fee00ff01100fe00ff001110e000f000122ff0000f1233e000ef0ef11f00fef0ef10000fe0ff010000ffff011000000000110000000100fff00001100f000ff00000ff010f10000ff010000000f0010011110f101001110de10100011fdf01100111edf11001110eef100011100000000011011110000111000010000000ff1100000fff0011f0100ff0f11010ff000001010010000000111100001001101100000011110000000000000000001000110ef000000110ff00000101100000110f02110011feff1210f01ffede1200010ffde11100100edf01111100ff00100110100000001100000000001100111f0022100f000001110fef1210110efef022022efee0f22031ef000022f420110f021f4200000011032ff000110f210fff0000000000000000010001110001100110000001111111010f012211111000000fe221100feff022011f10f00110100001001100000111011000111210100000000000000001011110001100000010000000000100000100101101000ff001111fff0f001011f011000100100011001001100100000f111010000000000000000001111122200110001002102110f00011012000fff110120000df0101f0110de110001222fe01f110111fe11011111100110111111f0100110000000000110f000000110ff001000100ff0011f0100ff0011f110ff010120100f0120121102eef00021022edfff011013fdee00100111fff011001110001000000f00fff000ff123edf001f1123fde012112121de114440001ef0032ddeefe2f11ed00ff2201fdd13011200eddf10001000fef01001000000000000000f021000100f03220ff00111111ff010122ff00f000011ff0ff000020dddf1000110eef230000f10f23ff00fe01120e0000ff0110f0100000000000000fff0fef0000ffef0eef0000f0120fe00101121100011002200100110f000011001111111000001220f0ff00feeeefff000fedef000000000000000000100fffef0f0100ff00ffe100100100f00001111100f0f0011320000000fe0201001ffedf10111fefed0111120fedd11102110fde0210112110010000100011fee000011210ff001132001f0101430f01001013feef0101f020fee0100f020fffef0100210feef0101111ffff100121200001001110000000000010f0000000010f1100000010f00000001100100010000000f0010f00f000101000f010000000ff0ff1100f000fe01101f010ff0100000000000000110010fff00000000ed001000fffedf02110f01ed01121ef01fd12f0ffffee122ff10fee0401e0100012101ff1001121010001112000000000000000000ffffeef00ffffffef0000000f01ff01010f021fff001ff1200ff0000131f101ff0110ff0110000ffff101010fe000000110f0000110011000010000011000110001100f000000110fff0010011ffef0010010ffff000112fff0000001111110001001001000110011000000000000f000000000000000000ffeff0221000feef011000ffef0111f000fff0010ee10f021f1ffe10f132f000d10d031100fe11de22100ff00dd12111ff00edf2101000000000000001101f0110001000f0210f01f000010f000f010010ff1ff1100100e1ee1100000e1ef0111000e1fe0210000e0ff0210000f000110f0000000000000000feee0001100eef000ef110ff000fdf211000d00de010fff010ff001102322220f0221f0321eef001010fddffef010fede00ffff00fff00fff00000000000000000000000000ff1101000000010010000000111110100001010110000010000000000100000f00001000000110010000f01000000000000000000000000000100000110f000000111000001101211011010fff11011fef0ff11011ff0110010100f011000000001100000001111000000000000000000f0100edf00f0f11fddd000ff20dddd011011ed242ff100014443000011f00d000ff0fffde000fe000ff0f000000f000f000000ff01000000010000000111001110011100010100000ff010000011ff00ef0f1100ffee0102001010111011111100110111100f010f01000f0000f011fff00000000000000000000000ff000011000ff000000000ff00f0000110e0000ff1013e01f0ff0f23f11f000ff22010f000ff11010000fff11100000ff011000000000100000110f000001210fff00001110ff0000011000f0100001011011010000111100100001111101f0000110111000110001000f001f0000f0000000000000ff001100f0ff011210f00ff001100011f10000001210100fff0f12110ff001e011210100000102111000000012100001010111112100000f0000000000000ff0100011100f0100110010001001101f0000101110ff0f010110ff00ff20110f010ff20110ef0f0010111ff0f01100110fff00000000000000000100fff0000000f0ff1100000f0ff2200000f0ee32f0f1000ed42f000001dd41f00f000ee41001f010f0110010010000001000f000f000000000000000000f00000100fe0fef00100feff0eff1000f1210ff111fef0023f110f0fdf33002220eef211f130ef010010fede0200000fedef1000000ff0000000012211011100220ff00f00111ff000f00010f0ff0000e01121ffe00ef1130eef01ef2220f0010e0012200000ef111210ff0ff01110fef000f0000ff0000001100ff000112100ff1ff1110e0ff1f020ffeff02f020fff1001012000210011021f11df211011020df11000011ed011000010ee1100000000000000ff000fff00f0011110e00f0011110f10f0110010011001110000111010f01001100010010010000000000100000ff01001ff00f0100000000000000000f0010ff00000001fde010000f1fdf00f010030d01100f004fd111f10ff1f2110f20f00f301000f00f02010000000110100000010000000000000000000000000000000110f010000110000100011010101000001001010110f000000001010101000100100110001001010000000101100000000000000000000f011000ff00f0210000000f121f00001ff24000001feef3ff0011eddf30f0020fde12000020ef0110f0011ff01000010fff00100000000000000000000000001110f0000001100f010f0000100000f00000021ff00000e121ff00f1fe1210ff0f1ff0220ff1f0fff210000000f0110f00000000000000000000000000110f0000001000000000000001001110000001001110000f00001000011110010000011111100111001000000010010f00000000000000fee0fff0000fff00000f0001100f01000111220131021ff001120f2fefff0f10e1fe0111020e1ee0111010f0fef011000f10fe02000000000010000000fffffef000fffff0ff000f00ef110001110f0200f0111fe02010f110e24200f100ff10f000000f10f0000000fff100ff100fef0000000000000000000111101110011f0011f1000f00000ef000011111ff010232ff00f0f042eddeef0ef0ddff0f10ffff1212211f0002112210fff0110110000ff000000000feeff00000ffffffffe000ff0ffeee10f0000fdef20f1211ed2011000112320110de3220f102fdd321fef01eeef0fedf00eff00eef000000000000000011111100f0100010000f001ffff001ff11ffef011001ff0ef111010f1311102101110e011101221fef1110120fee01100210fef010000000000000001000f00000100000f00000111210110001112102100010fffe110000ffeef11011f00f0110100010f11111000000100100000100000000100000000010000fee0000f00ffe010f1010f0232101011244211f000100eef1ff0ffeed00ff0f000f00fff00000eff0f01010ee0f0f111100ff000001100000000011000111001100001100000011011000f0110011011f01ff0f1011000fff011011fff001110000f0100110000010001100001000010000000000000011100000101210ff000001100000ff0000001ff0f00ff110ff0010e0010ff0000f01110f0010f011221001000111110000f0010000f000000000000000000010000001001000000000000000000000011110000f000101010000100011000110100000011000000000100100000001101100000000000000000000f0fff01000ff0fff00010f0000f00000e0101ff100ef00f4ef1f0f01f14e00ff000e13e0fff00ff21f00000f001ff00110f010f000000000000000011110010f0112100110f10020eff00ff011fe0010e0110000110efff002111000ff031fff1101121fe000012220df00001111fdf10001110000000000100000f001100000000000000000000000000101000f0000101101000101011010011010100111100100000110000000f110001100000000000000000001001000ede02200f00ee01231ff10ef22111f011f03200fff00000e000eef0ff21133ee00df321220e00de13221000fdd010f00000fff00000000111000111001111f0001001110eff0200011fdfe0100021fede0000000eef1110000210021ff00122f110f00122111fff00010110fff0000f0000000000000f0110000100001101111000e0000100f00e000000ffffe0f000fee0edf0000f0ff01110f0001133110ff0001110f00f000100ff0000000000000ffef0100000ffe010ef200fff011ef1010f1012df2110fff0fd02110fffffd01001122232100ff1101430f0eeff0231fe0fff00120ef00ffff000f000000ff00000110fe000000100fff00000111fef0111f10000001110000132100100000001101f0000ff100f000100011ff0f010f010ff000000000000000000f021000110fde00001000fdd0f0f2100eddef1122feede121021f0e24221110de0411201120e22efff0031f20eef00e00010ff00000000000000111110111000100010010000000000100f00100001100110fff0010000fff0100010010000000100000001001001000110001000000000000000000000f0011000000101110001000011010010001110000101101200f011100f000001010010000000100110000101001000110001000011000000000000000000ff0110000000ef010010000ff000110ff11fff0000f1320f10000133210110100f010010110ff10f010010fef00000010fef001000000000000000110ff000000000ff00000000ff0110f0000000110f0ff0000021000f001ff2200f000fef211001000ef11100100ff001010100ff00000011000000000fefffff000fff00000e0ffff11111f0feef1122200eee001211fffef000001ff00ef1ff110f1fde20f02002fdd01001002fef0000100000000111000011000110001100f0100000000f0000f0000f00011f100ff011210100ff112110100ffe01110110fff01110011fef001000110ef1110000000000000011000ff000010ff000001010fef00f0100feeffee01ffee132fe010f02311100101332f0100101231f11000f0010f000f00fee0fffff000f00000f0000000001110f0000f01100f000fff1110f0010f02100011fffe3100010eedf2000010ddd01100011ee0100000120e0000001110f000000001000000000fff0ff00000ff000ff100001100000000111120f00000ff021f00000edf21000000fd132101000fdef01000000fef00000010fef0000000100000000000ff0011000000f000111011feef022000fedeff11100ed010000100ff3123ff000122e1300f01231e01ff00111f000fe0000ef010ff00fff00000000ffeff001100feff0ff0010ff001ff100000001fe101110101ff100111100001000000f0101000ff001111f0fff000100f00ffff0000f000f00000000000000000f00000f0221f0ff0fe01220ff00ffff041000f0f0f032110fff1f001111f00ff1f0111110f0fff00110ff00f0001100000000000000000000011000111001110ff00100010ffff1100000ffff110010fffe011011fff0010001100001000011100001000011000100000110f010f0000000000000000fff00ff000f00011fe00000f0120e0000000122ef00ffef143d00fffef143e010effe121e01ff0ff010f010f0ff110f01fff0021000000000110000000ff0000000fff01220f11fe0121100111f100111011001f00f20100000ffe101fe01000f0f1fe00000f0f0001100ff00001000f00000000000000000ffff011100ffff1ff0210f00011d00000f0f01e01110f0f0fdf1010eff10f01f0001114420ff0111134fefef0110fedd0ff00ff0fee00fff00000000fffff010000edde002100fdde0f01221edf30f10221ef12e0314ffe10fe240fee130dfe22dee130eee0eeef0110fffeff0001000000000f00000000000000f010000f000ff001000f0fe000101101ef0000f2010eff201f21220dd400f11120de20101200dd11000111fdd22100011edd120000100ff00000000000f011000000ff010000f00f0110000f0011100f10012211f001001111100f00fff01000f00fef00000f000ff0001000000ff00100000000000000011000110001100ff00100110ff000101110f0f0010000000000100000120000010f00100f00100f0000f0000100000000011000f00000000000000000000011100000000111100f000f001000000ff01100000ffff11f010ffde011f0110fef11100110f01110f0011000000000000001000000000000000;
  initial weights_NN1_layer1 = 48400'h111f00fddf01ff000ffee0fdeff21ffd0fdef141efd1ede1343f0e0fdf024211e0feff33f10ff2edd43011003ddd01f0f101edeffdf110011000f0000000f0ff11000ffffee00f00ffffedf0f011100edff00010111f010f0000122101f00ee3201f0f02ed1331dff01fdeffedf0000ffffef0000000000000010010fdd00110fffee01f01fdeeee00ff1fd021221fefde204421000f22dddee0f0331edefe0f0121d011001ff10df100000f00ef0f000000000000001100ed02201210fede111122211ee111112232fd100111233201f00f13210f1ff0df10ff00000ff00ff01200ff01f001100ff0f0f01000001110000000edeeee0000eddf21f0f00ddef3201f12fff131f0f12fe121001e0111330e01df0f23ff100effdeee232fe0fdddf221ff00dddf0100f00fff01100000000000fff0000000000ff000001121000f0110211110001f0fe21110ffe0ff21121f00001111100000000010000010000000111000000000000000000100000fef0f00f0fffffff00f0122ffff001111310f0010fff131f011edede330001ff0dd231000010dd23111001ddf120110ffdef0100110000000000fff0ede000ffefeddef011feee1f0f0210ef4430ff100f24411f0f01121f01f0f0121ff0f0ff001ff0000f0ffeee101000fedef00110011000001000fff00feff00eef0211100fedf11000000ddff00f000100e0220ff011f032e010011134fd020f01232de1fff0101ed01ff0120fed00f000000000000000feffedf000ede1100ff00ed134310e0fde034420effef2332f0e0fe120fd00d0fdeffdf20e01ddf10110001ddf221f1001ddf110010000000101100011100fef11010111fdd11fff0120dd3100f1110df42ff0f000df310f100ffe01000100001100f00010000000001000000001110010ff00010000ff0000111112320f1210110021f10120ff011ff0120f001011100fff011210ffee0010120010200001100122112001101121220f1210210210000f0000000000f100f0000ff122fef00111211fdf011101010fe01232fef1000122ddff0030010dffee14000edf0002200feff001111000ff01210000000000000000100112210f00000100000f0000f01000f0010f01111ff001f11011010fe0101101000f00011010ff012110020fff21110010ff02000000fff0000000010ff022100221fee121f0321fde02201320dde0031230deeff02134eef22f0313401110f021232000ff010222ff0f01100210fef0100001100000000010000110001000010100000001001100ff0100002010011fff0201100ffff11001f10ff111001000001110010010101000000001000000ff000000000210221ef1ff00112fde1ff002010de0ef10ef1fde0de201021de1ee43330eef3dd4200dee23e031ffdff12e021eeef0120000ffff011000000000000f01111221000111000f210110fffff11010fffdff2101100f0ff210200443e0110111241ef111110121ff110110000ff010110000f000000000000000010001110001111111000000111011000e0121101211f0000fe211200efff021121f000011111000000011000011010120001010101100000001010000110f02100011feef1110f00fde114000f10ee210e020eeeedddd02100efff11f3333203443f0231002120fff0eef100f0ff0fd0100e000ff00000000000ff01100f010f01420ff0fee01341ef000fef142ff101fe01340100ed100f1121fd1e01e11221fff0ef001230efff00002210000000000100011000f0111ff000ff111ffff110000010fff1101010edf120112112fe020012443fef3000243eff020f021ee1011f0110fe011102110ee0100011100011000fff0022f00000f0121e000fef0020d000f011f31df10100ff22d1102120d12e0001220d01000020fde000100110de00110001fde011000000000000000001fee010001221ddf11011023ed0210100221d112121f000e011010efe1300001fdf120f1f001ee00ef0f0010f0ffff0000001000000000000000000110ef01000000fee020f00010ff110f11110101ff010f20f11f2000122102111000f0fd01100110fddf0000031edd00000122fde00000011000000000000111100ff121001010ff110ee0000fff1efee110feeee01121100ddf22210012dd12f0000221420f000012320fffff002210f0f00001000000000000000fedf00f0220fddd0000220ddddf000110edddd0f1200241dd0f0103442ef0fed0f02f210fdfffff1210fffffff1200eeffe01110000000111000100110222000e0112111f1ef0132001f0ef1210111f1f0220ff1fffff0f0010ee0fe11133fed0ef0f2330feff012331feeff021210ff000ff00ff00001000ff000000000f021f0000011011000f0120e11ff1f0210e02fe10e120d12fe10d03fe21ee1edf3fd32ff0fe02ff110f0ff01ff100000110000000010001fdde01002221fee100134222ff1f0343001001f032ede1101ff100def0f1ff120efef01fe023fffd110f03320ed10011131ff0100111000000000f0000eee0100000000e000000111ff00112111111101121101211f110010111101202101001f0101100001000000f00000f010f01f00000000000000fef0f00ff00eff0fff001fff01f10f00f0000120f0002fff14001001fdd442010f21dd023000f13fddf00f0ff22dd00ff00122fde00000011000000000220f021100121ff011f01000ff011ff10ffef011fe1fffef033ff100fff2430f00f00e1320001ff0f03200111fff221f0011fef220000000000100000010fffef000111feeddf01000feddde1100ffe010e0000f02312000011031f320f0eef2dd32110fe20de22001102ddf1110ff0fdf11000000000100011200110001210f011000100f0010ff000ff0f01f0000000ff1e0100111edfe11e12221ef021ef012222120ef101212100ef000111ff00000000ff00011110000f0122100011f011100010f0000011f01f1111120f0100001000fee0100f0011df0100f00111112000001101110ff1110f100001110000000000010001100f1211ef10001011ede0f001110eddff1022eeede11f031e213312122fd022e02032fd040df10110ef2eef1000fe00ef11000000000000000111100f0f01111100f0f011ffff001ff110fef012000f00ff112011f0200102013111df11201211fdf11101100ed021101100ee010000110000000000ffffef00111fef1f001111fe12ff01210ff11ff01000011fefe0000033ff0f00003300000000f22000f000ff0110ff0000fe010f000000000ff00000fef0ff0000fef110ef020f0011fede201fe00edde1f0ff0000011f1132114210f120f01eeffff01220edd0fef0210eef00eef10fff00000000000000000000000000001111000010111110010f0132000011001220f10000110f0010000110f00001000f0100010010110f01101f011f00110000000000000feeff012100efeff021000ffef01210f0fff00222ff1ff022200ee1fe013101ee10df210120f00eef10020f01fde0f120010fee001100011011111000feefff0f000eff00010f0ff010012100eff01122200fff0014220f00fff2201ff10ed00ff0ff10edefff000110ddff0100111fff00100111111110000112110110001111f0111001010ef100000120e01e10f0120effe10f100fe0011001011110f00011121fff00001110f0010f01100f0000000000000000000021eee000100110ff00f000010f01f0010011112f0010002202f210f201102022222f10f2f121001100100100001001f0111011f0000f00f0000000001100ff0fff120000f0fff0fff01f00ff000011f0100001f21f00010edd41f0001fedd11f0000feef120000feff0110010000f001000000000000000ffff010000eeeeef2000edddedf2210dddeee01200ee1411002ee02222420ffe23002220fee22eef1100ee21feefefee010f000fff000f0000000000000000fff010ff0000ff00fdeeeeefee00ddf21ffde00e1423200ef01311231feffe0fe210feefe10121eef0ee0210fff00eef000fff0000000000000000ff00ff01000e0110ef0010ef121ff110f00212fe10ffff033fe20efff1430f1101fd032001000dd130f0100eef21ef0000ff031f000000f011000000fef01110110ff00001011f01110120221fef10120332eeeeff20231effeef30340e000f02124fdfff0121230feef1310110eeef2200010100011000f0000010000fffff0111f00ff0f000ff1100e0f00fd2000ff0101f200221e310011121dd21101221dde1210022fdd02200021eddf11000010ff0000000f001100f000011110ff0f0001100001ff0111111110000f111101100ff01110101211010001011101100010010010001100011010000000000000000000210001f00f020ff01e0fe02fdff0e0fe1110433feef12143f10fe0f1ffddd0fd1212edddffe1103feffffe1221fef0f0ff121ef000000000f000000edf00f0010ede021fd021ff1211fe122f03101fff24232f00f0e0221eddf1fef0e02f022fdfee0322210dfede232210f00ef021011000fff0011000000ff0022100ffff1001111ffff0fe00110fff00e00010ff021e0ff00f0010ef0ff001024100ff01001230ffff00f1220e0fffff010ff00fff000ff000001200220f00ef0e0210e00fff0120de1ff121341ee0ff10e030eeffefef13fed0ff00132fed0fef0221feefee01220fff0ff011000f00fff00000000110fedde0111ffe0dd011100ff0fd1111fff021d0311110010d2410f1100dd4211200ffef41102f01f0121001000f111000100e011f00001000000000122110000002221f011100220ddef000011ddeef0f0f00eff01001f0122fe0111ff22fed0101f0210ee1101f0220f0100000111000f00011000000000000f00fef010fef00fde020ff110fde01001210fef1f03320ff101ef440ed0202ed3eddd1212dfddeff0101fefef0111210eff00111100fff000000000110000000011100fff0000100000000ff0100100020010ef0f111110efff010111ff211110100001111101001f010100101100100000000000000000011100f010001100fe0000121ff0ef000022f0fe0110f1111ff121002033001120020fedf0220030fddf0110120eddf0011220fdd0100012210010000110f01eff0110ff23fef11f0ff1110f10ee011010110ee011ff0010ff11fef00100143e02201ff142f121f1fff111310f1ffff2231ff00feef1100000ff00f02210f0010ff2200fff01ef220ffff00f01100010fe00210010fdde142f0110eef132f0111fd0011f0013feff02000111ff01100001100111000000ff011001120f0f01f12120f000101121ff011001110003110010101430000100f1101101110f01f00011011000111f0f11001110000001111000000100ff02101100fff020f0f00f0f130f0ef100023ff1f010ff03ef100f0fe030e10ef110020f1fef111220f000f111000f00000110000000000000000fee0f0110000f010121f0120f00011f010f0210230f20ff00013fe2feeffe020d20de122020d2ede222020e10de131110f10ee121010000001111000001111ee00000110ede001ff221fde111ee0342ef101ed0432ef1f0ed0002000ffef0013100ffe0ff01000ff0011021eef0001222fef00011000ff0000f000fe0210f0001fe020100f011f120110e0100100021000111ff022010f20fff101fdf3000f0f0dd02121f0ffed0112001feeef1110000000100000011100000f0110100111f00f00f111200fef01fe0221ff021fdd32000110ede11110120ff21210f22100012100121fff0100ff11ff0f0000f0000000000012211110ff02320ff110100100ff10121fe10011011110110fef112f0eeeddfe0fedd01ef0f10e02420110002221111000012100110000000000000fef22111001f0312100102123f00ffe0232fe11def022ede01ddf020edeeddf1100011e13210ff112343000fe0023310f00ff01320000000000000000fff00011000ff000121f0000100022f0ff000f0130000fff0103f010feef1120011fde02111010ffe0001001110ff000001f0000100000000011100000f01000000f01111000100100110001101000100f00110f121ff10200f1100010100f1020f000000110e000000011f0000000000f010000010000000001112110f00121100000000110ffff110121efeff22f23ffff0f12f23ee010f12e341010ff12d340f10ff11e23fe0f0111f12110e0010011100000000010ff0eee00011ef0ffe0ff10d0121ff000fef104df0ffed1e14df0ffdf1d34d01ee11fd23d1fff00ff20f1000fff00ff00110ef00f000000000000000110ee0f00011ffeef000020ff11ff1f02ffe01002ef00f022e02ff0ed243df1e12fdf43f01e131dd21102f020dd002010121edeff01000100ffff0000000f000000110f0ffff1011000ffff0f0010011100010f0022001011f01110100111311f110f0111101110f1100101100f0110110f0000f0000ff000000010f000000fef0ef21011fde0ef41010edd0df4100fee01de2111ee234201011342e132fff033fd01edfef0eeffeed0f00de00ffe000ff000f00001000010000f2200e0f000f212fee01200210ff12220021dffe3200030dddd1300030dddd122103fdde11120242ed000110223ff001210011100011000101111011011100110120120f000f02111000000f21011110eee2111f111eef1110e120f0e100112221fe000111220fe10f12110ff01000000ff00000122131fde002322100ff101421f00f02e032fee0f12e042eed0003ef41fddff12e0420fef003e04230efef200222feef11012230eef000111000000000000f011100000000222f01f0101222010000000f111ff11f0fd011ef1000ef001fff112f00f10ee020e00f010011ff00f111110ff000000000000000fddde01210fdddd011101fdffe000000001000ffff0110032f00e020f1442220010e0322110f20de12101ff10fdd0f00f000edd00f00000ff0000000000000f022000ff0ffe11101011ffe010f00110fefe0ff00fffef00f0f0eee132f0000f13320f0001211eedf001220feee00f1110ffff000000000000000000fef00f00f00eef00e00f10f0000eff01101210e0ef0020210110021dd10f100020dd20000e02dd022001f1fdd01201100fdff000000000000000002231ff00ef003200f01fff02210de1ef00220ede1e022310edf2d012410de02d01f130ee01ff01100ff11ee0220df011fef12fde0000000000f0000000001000000000110000000011000000f0012100101ff0110011100f00f0011100010f1100000010010000000000100000000001100000f0000000000fffff01100fef0feef100ff010eef0010012fef01001111f0122ff0f1fe2301f0ff1023ddff10e123edeef10ff1fffff00ffff10f0000000000000000000ffeef00100feefff01121ff00f011021f12fe111f11122f022fff2131e312ef11f0dd211f01000de1111110f0ef00012100ee00000122100100000f00ffddf000ffffeef0011000ff23301011f0344410f000240f22000001eddf100f0f0ee0eff0ff0fe00ef10000ee21e00110ff010000000000000000010ffff0001110fe010001100f0110000000f110200ff001110200f0ff11f031001fef0f021011fffef1210010ffe011000110ef10000011100000000000110100001001101110100110ff110001320ff101111330001001111ff011000110000010010011101100101100121000000001100000000000000000010111000000111220ffff012110000ff021fef00f001ddde000f0ff01110000ef210110012122000ff001221000ff001100100ff000ff000000000ffee122000fedef1341f0effffd240e1010efe13fe0ef0f0f23dd10f002242dd2ff12023ddd0123001fddff111110ede0fe0f010fff00dde000000000000ff1100f0f00ff110001010e021f00112fe13100011edfe30e1011ddd240e1031ddd23f01122fd040e000120d140f00100fe0110000000f000000000000ff00000010fef10f0ff0fee01ef0feddfe01eeffee221120f0f143114100f0230df0f00f0131e0fe0000010f0fff000f0ff0fff00000000000000110f011201220df0ff11221fd010e11121ee0fff00002132ed001f00344ee0f10ef3320fef1fff24310df0ef01221fde0ef11131edf000f000fef0001110f01000120fff000f01000011fef001f00f01f0010f00ff0f1100010fedd10f12212f0020ef012233110ff00211100feef0f010ef000ff000ff001000feffef01100feefee01010ff02edf10000f140ef10fff02112f1fefe10d4300001f0ef321ff1000e11000f000001f000ff00f00f000000000000000001002210f0ef21f201000ef1021ee012000123def00021011def00111d0fdfff11dd141dff000d2411000fff021e11000ef010e010000f00000000;
  
  reg [(hidden_layer*out_layer*weight_bit)-1:0] weights_NN1_layer2;
  // initial weights_NN1_layer2 = 1200'h1fe1f0dfe02ed112d0f002f10fd2101ef0ddff0ddeee1e111021020effd012200f01f1e2100f22ff1fdf0fd2001ee2f0ee1000020ff10f01f1f10e1d02120d2e2fee03f1fe01ef0012f2ef0021f0f2e0fe0ed2f1f1e021dfee0efefeff1211fffe020fe0df022f10f0df0d1010e01f2e0d011f20f1f1110eeff23f12fe10f1f12edd1f1ff00fe1ff10f0f0e1ff102fef1102ef0e0f1e;
  // (200 Neuron Attempt) initial weights_NN1_layer2 = 8000'hef0010f0ff100020f1000000f0f010001ff00e0f10f00e00f0f00000fe0f0f0f00100fe010000f0f000000f00f0000000e0f11e11010f111f000000e01f01f00e01f0f1011f00000ff00000000010e0001f1f0f0000e000f01f00000f0f1001f1001e0ff0ee00000f010000000010f000000d000ef0000f000f00e100000000f0000000f000e00f00e00d0000000f00f000000100f111ff1f00f000f0000f0111ff0f0000fdf0fe0f0000100000010010f000f01000e0ff000001ef001e0100e0ff0100000110000010000001f101000000f00100010ff0110f0f1f0000001f0000f010f10000fff000001f00f000001000000000f00f001f000003ef00100f0f0000001000f0f0f0f21000000ff0f0f1f0f0f10ef0001f00f001000f00001000f000010000f100000ff10f0000001001f0f0e00f0f00fff000f000f000f000000000111f000fff0f01f0010000f000000f0f01f0fff00e000000f0100010f00100e0020000ff000000000000e000f00100ff10f00000f0000011ff0011100f00000000000100ff0f0000000ff11ff00100000fff0101fe00f000ff0000010011f0000f0f000001000000011f03ff11f0e020001ef0011f00001f010000020ff00f00f0120ff002f000001010f00f0000010fff00f001000e00101200e0101101f0001f000100f0100000f0f0f01000000011f001000f010fff000010000001f001f1f0e10f10010fff00000f00001fff1f10002000000000f00000f000000000f00e0000f00f100000fff0000010f010ff00e000f001f10f001010020f000ee000f0f000010f01010e00011f00000f0f0f000efe00ff00f0ff00010101010100ff00101000010f0ff0f00f01f0001ff000000010ff101f0f00000100f001f1000ff00000000100f00ff0f00f1f100ee00010000f000f000f0010000f0010e0010100000f110001010e10010f0100fffe01000000e00ef0f00e1000001200000f0e01f10010011100001f000000f00f010000ff0f1000f00010000000000000001100000000f10000000000101000000f01100f0000f0000e00011f0ffff0f00f00f0f000000000100000000f00f00000001000ff0f0000f000f1f0001fe200000ff0f100f10000ffff100000f0000001f0000f011fff0f01f00f1001001f102f1f0f0000f01f0f0f0ffff00f00f00000000000010000f000000f000f00fffff000000ff0101010f10f00ff000f0f00ff101001ff0000ff0f12ff10f00000000000000000010000f1000ff00000e0f00000ff000ff0f00100000010000f00000001000f00000000f0f0f0f000f0000ff00e0f00000f0f0000001f000f00f000ffff0010000001000100e0ff0f010100100000ff0000f0000000000001f000f000f0f00000011ff00;
  initial weights_NN1_layer2 = 4000'h110010f0ff0f10e0fe0d0effff0001110f01ff1f000f0f210fd0e1001000f1f0000f1e000f010fe00f0ffd001f0001e0001edfe010f01e00e100f000000e020ffe100f10d00f0ff01f0f0f00ee0f0e00000100e100f00f1011d0d01fd01f001111e011100f100010200f10e0f000f1000010100f0ff0f1f0100f01100f10f101100f000f00f011110e0e0f1ef000200000000021df0200f000f0001000001000f011f0fef01fff0000010ff0100efff0f1fe1020f0f0fe1f011000fe11000f010001fff0f1ff00f1f101e0fdfe20100010f100221fd01e020f1000fffff000100100100120f00f001010001f001110fff0010000fe00f2010101101100f110f0f0e0e002eff00ff10100e0010e0100f00f11eff01000e0fffff00000010f0fd10ff000110002f1f11ff000f000e0e00f0fff0f00f00f00000f1f101102f0100f01000f1e00000fef0fe00f000100f00011100d00f10f1f010210fe1eff001f00f0111ffff00000f1001f0111101e1101000f0ee010d011100e0000100ff00f211fdf0000010010df010f00001f010000f12f0ff01f0f0fff01e0f000011ffff001ff2001f00f00111f1f1f0f101f1ff0fff0ffff0f01f1fff010100011ff00010fffff0ef010ff000010ff001ffff0f0f01f0f000f0f0f00110001f110f101f0f00fff0e0010001e000001f0ff00ef0001ffe010;
  
  integer clk_counter = 0;
  integer clk_counter1 = 0;
  integer clk_counter2 = 0;
  wire clk3;
  wire [(hidden_layer*4)-1:0] hidden_layer_out; //30 hidden layer output with 3 bits each.
  wire [8-1:0] output_layer_out[out_layer-1:0];    //10 output layer with 4 bits each.
  wire [output_bit-1:0] out;
  //assign clk3 = (clk && !(clk_counter==0));
  reg [8-1:0] max;
  wire [WIDTH-1:0] div_num = 6'b000101;
  
//integer i;
input_reg S0(.reset(reset2), .clk(clk3),.input_features_in(input_features0),.input_features_out(input_features));

always @(posedge clk3)
begin
    if (reset2)
    begin
        clk_counter <= 0;
    end
    else if (clk_counter < 3)
    begin    
        clk_counter <= clk_counter +1;
    end
    else if (clk_counter == 3)
    begin 
        final_output1 <= final_output;       
        clk_counter <= clk_counter +1;
    end
   
end


always @(posedge clk3)
begin
    if (BTNR)
    begin
        clk_counter1 <= 0;
    end
    else if (clk_counter1 < 3)
    begin    
        clk_counter1 <= clk_counter1 +1;
    end
    else if (clk_counter1 == 3)
    begin      
        clk_counter1 <= clk_counter1 +1;
    end
   
end

//Neuron_NN1_layer1 N1 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[483:0]),.bias(3'b000),.out(hidden_layer_out[3:0]));
//Neuron_NN1_layer1 N2 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[967:484]),.bias(3'b000),.out(hidden_layer_out[7:4]));
//Neuron_NN1_layer1 N3 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[1451:968]),.bias(3'b000),.out(hidden_layer_out[11:8]));
//Neuron_NN1_layer1 N4 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[1935:1452]),.bias(3'b000),.out(hidden_layer_out[15:12]));
//Neuron_NN1_layer1 N5 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[2419:1936]),.bias(3'b000),.out(hidden_layer_out[19:16]));
//Neuron_NN1_layer1 N6 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[2903:2420]),.bias(3'b000),.out(hidden_layer_out[23:20]));
//Neuron_NN1_layer1 N7 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[3387:2904]),.bias(3'b000),.out(hidden_layer_out[27:24]));
//Neuron_NN1_layer1 N8 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[3871:3388]),.bias(3'b000),.out(hidden_layer_out[31:28]));
//Neuron_NN1_layer1 N9 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[4355:3872]),.bias(3'b000),.out(hidden_layer_out[35:32]));
//Neuron_NN1_layer1 N10 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[4839:4356]),.bias(3'b000),.out(hidden_layer_out[39:36]));
//Neuron_NN1_layer1 N11 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[5323:4840]),.bias(3'b000),.out(hidden_layer_out[43:40]));
//Neuron_NN1_layer1 N12 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[5807:5324]),.bias(3'b000),.out(hidden_layer_out[47:44]));
//Neuron_NN1_layer1 N13 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[6291:5808]),.bias(3'b000),.out(hidden_layer_out[51:48]));
//Neuron_NN1_layer1 N14 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[6775:6292]),.bias(3'b000),.out(hidden_layer_out[55:52]));
//Neuron_NN1_layer1 N15 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[7259:6776]),.bias(3'b000),.out(hidden_layer_out[59:56]));
//Neuron_NN1_layer1 N16 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[7743:7260]),.bias(3'b000),.out(hidden_layer_out[63:60]));
//Neuron_NN1_layer1 N17 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[8227:7744]),.bias(3'b000),.out(hidden_layer_out[67:64]));
//Neuron_NN1_layer1 N18 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[8711:8228]),.bias(3'b000),.out(hidden_layer_out[71:68]));
//Neuron_NN1_layer1 N19 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[9195:8712]),.bias(3'b000),.out(hidden_layer_out[75:72]));
//Neuron_NN1_layer1 N20 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[9679:9196]),.bias(3'b000),.out(hidden_layer_out[79:76]));
//Neuron_NN1_layer1 N21 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[10163:9680]),.bias(3'b000),.out(hidden_layer_out[83:80]));
//Neuron_NN1_layer1 N22 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[10647:10164]),.bias(3'b000),.out(hidden_layer_out[87:84]));
//Neuron_NN1_layer1 N23 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[11131:10648]),.bias(3'b000),.out(hidden_layer_out[91:88]));
//Neuron_NN1_layer1 N24 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[11615:11132]),.bias(3'b000),.out(hidden_layer_out[95:92]));
//Neuron_NN1_layer1 N25 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[12099:11616]),.bias(3'b000),.out(hidden_layer_out[99:96]));
//Neuron_NN1_layer1 N26 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[12583:12100]),.bias(3'b000),.out(hidden_layer_out[103:100]));
//Neuron_NN1_layer1 N27 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[13067:12584]),.bias(3'b000),.out(hidden_layer_out[107:104]));
//Neuron_NN1_layer1 N28 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[13551:13068]),.bias(3'b000),.out(hidden_layer_out[111:108]));
//Neuron_NN1_layer1 N29 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[14035:13552]),.bias(3'b000),.out(hidden_layer_out[115:112]));
//Neuron_NN1_layer1 N30 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[14519:14036]),.bias(3'b000),.out(hidden_layer_out[119:116]));
//Neuron_NN1_layer1 N31 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[15003:14520]),.bias(3'b000),.out(hidden_layer_out[123:120]));
//Neuron_NN1_layer1 N32 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[15487:15004]),.bias(3'b000),.out(hidden_layer_out[127:124]));
//Neuron_NN1_layer1 N33 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[15971:15488]),.bias(3'b000),.out(hidden_layer_out[131:128]));
//Neuron_NN1_layer1 N34 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[16455:15972]),.bias(3'b000),.out(hidden_layer_out[135:132]));
//Neuron_NN1_layer1 N35 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[16939:16456]),.bias(3'b000),.out(hidden_layer_out[139:136]));
//Neuron_NN1_layer1 N36 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[17423:16940]),.bias(3'b000),.out(hidden_layer_out[143:140]));
//Neuron_NN1_layer1 N37 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[17907:17424]),.bias(3'b000),.out(hidden_layer_out[147:144]));
//Neuron_NN1_layer1 N38 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[18391:17908]),.bias(3'b000),.out(hidden_layer_out[151:148]));
//Neuron_NN1_layer1 N39 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[18875:18392]),.bias(3'b000),.out(hidden_layer_out[155:152]));
//Neuron_NN1_layer1 N40 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[19359:18876]),.bias(3'b000),.out(hidden_layer_out[159:156]));
//Neuron_NN1_layer1 N41 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[19843:19360]),.bias(3'b000),.out(hidden_layer_out[163:160]));
//Neuron_NN1_layer1 N42 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[20327:19844]),.bias(3'b000),.out(hidden_layer_out[167:164]));
//Neuron_NN1_layer1 N43 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[20811:20328]),.bias(3'b000),.out(hidden_layer_out[171:168]));
//Neuron_NN1_layer1 N44 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[21295:20812]),.bias(3'b000),.out(hidden_layer_out[175:172]));
//Neuron_NN1_layer1 N45 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[21779:21296]),.bias(3'b000),.out(hidden_layer_out[179:176]));
//Neuron_NN1_layer1 N46 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[22263:21780]),.bias(3'b000),.out(hidden_layer_out[183:180]));
//Neuron_NN1_layer1 N47 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[22747:22264]),.bias(3'b000),.out(hidden_layer_out[187:184]));
//Neuron_NN1_layer1 N48 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[23231:22748]),.bias(3'b000),.out(hidden_layer_out[191:188]));
//Neuron_NN1_layer1 N49 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[23715:23232]),.bias(3'b000),.out(hidden_layer_out[195:192]));
//Neuron_NN1_layer1 N50 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[24199:23716]),.bias(3'b000),.out(hidden_layer_out[199:196]));
//Neuron_NN1_layer1 N51 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[24683:24200]),.bias(3'b000),.out(hidden_layer_out[203:200]));
//Neuron_NN1_layer1 N52 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[25167:24684]),.bias(3'b000),.out(hidden_layer_out[207:204]));
//Neuron_NN1_layer1 N53 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[25651:25168]),.bias(3'b000),.out(hidden_layer_out[211:208]));
//Neuron_NN1_layer1 N54 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[26135:25652]),.bias(3'b000),.out(hidden_layer_out[215:212]));
//Neuron_NN1_layer1 N55 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[26619:26136]),.bias(3'b000),.out(hidden_layer_out[219:216]));
//Neuron_NN1_layer1 N56 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[27103:26620]),.bias(3'b000),.out(hidden_layer_out[223:220]));
//Neuron_NN1_layer1 N57 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[27587:27104]),.bias(3'b000),.out(hidden_layer_out[227:224]));
//Neuron_NN1_layer1 N58 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[28071:27588]),.bias(3'b000),.out(hidden_layer_out[231:228]));
//Neuron_NN1_layer1 N59 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[28555:28072]),.bias(3'b000),.out(hidden_layer_out[235:232]));
//Neuron_NN1_layer1 N60 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[29039:28556]),.bias(3'b000),.out(hidden_layer_out[239:236]));
//Neuron_NN1_layer1 N61 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[29523:29040]),.bias(3'b000),.out(hidden_layer_out[243:240]));
//Neuron_NN1_layer1 N62 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[30007:29524]),.bias(3'b000),.out(hidden_layer_out[247:244]));
//Neuron_NN1_layer1 N63 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[30491:30008]),.bias(3'b000),.out(hidden_layer_out[251:248]));
//Neuron_NN1_layer1 N64 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[30975:30492]),.bias(3'b000),.out(hidden_layer_out[255:252]));
//Neuron_NN1_layer1 N65 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[31459:30976]),.bias(3'b000),.out(hidden_layer_out[259:256]));
//Neuron_NN1_layer1 N66 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[31943:31460]),.bias(3'b000),.out(hidden_layer_out[263:260]));
//Neuron_NN1_layer1 N67 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[32427:31944]),.bias(3'b000),.out(hidden_layer_out[267:264]));
//Neuron_NN1_layer1 N68 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[32911:32428]),.bias(3'b000),.out(hidden_layer_out[271:268]));
//Neuron_NN1_layer1 N69 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[33395:32912]),.bias(3'b000),.out(hidden_layer_out[275:272]));
//Neuron_NN1_layer1 N70 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[33879:33396]),.bias(3'b000),.out(hidden_layer_out[279:276]));
//Neuron_NN1_layer1 N71 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[34363:33880]),.bias(3'b000),.out(hidden_layer_out[283:280]));
//Neuron_NN1_layer1 N72 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[34847:34364]),.bias(3'b000),.out(hidden_layer_out[287:284]));
//Neuron_NN1_layer1 N73 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[35331:34848]),.bias(3'b000),.out(hidden_layer_out[291:288]));
//Neuron_NN1_layer1 N74 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[35815:35332]),.bias(3'b000),.out(hidden_layer_out[295:292]));
//Neuron_NN1_layer1 N75 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[36299:35816]),.bias(3'b000),.out(hidden_layer_out[299:296]));
//Neuron_NN1_layer1 N76 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[36783:36300]),.bias(3'b000),.out(hidden_layer_out[303:300]));
//Neuron_NN1_layer1 N77 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[37267:36784]),.bias(3'b000),.out(hidden_layer_out[307:304]));
//Neuron_NN1_layer1 N78 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[37751:37268]),.bias(3'b000),.out(hidden_layer_out[311:308]));
//Neuron_NN1_layer1 N79 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[38235:37752]),.bias(3'b000),.out(hidden_layer_out[315:312]));
//Neuron_NN1_layer1 N80 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[38719:38236]),.bias(3'b000),.out(hidden_layer_out[319:316]));
//Neuron_NN1_layer1 N81 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[39203:38720]),.bias(3'b000),.out(hidden_layer_out[323:320]));
//Neuron_NN1_layer1 N82 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[39687:39204]),.bias(3'b000),.out(hidden_layer_out[327:324]));
//Neuron_NN1_layer1 N83 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[40171:39688]),.bias(3'b000),.out(hidden_layer_out[331:328]));
//Neuron_NN1_layer1 N84 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[40655:40172]),.bias(3'b000),.out(hidden_layer_out[335:332]));
//Neuron_NN1_layer1 N85 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[41139:40656]),.bias(3'b000),.out(hidden_layer_out[339:336]));
//Neuron_NN1_layer1 N86 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[41623:41140]),.bias(3'b000),.out(hidden_layer_out[343:340]));
//Neuron_NN1_layer1 N87 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[42107:41624]),.bias(3'b000),.out(hidden_layer_out[347:344]));
//Neuron_NN1_layer1 N88 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[42591:42108]),.bias(3'b000),.out(hidden_layer_out[351:348]));
//Neuron_NN1_layer1 N89 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[43075:42592]),.bias(3'b000),.out(hidden_layer_out[355:352]));
//Neuron_NN1_layer1 N90 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[43559:43076]),.bias(3'b000),.out(hidden_layer_out[359:356]));
//Neuron_NN1_layer1 N91 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[44043:43560]),.bias(3'b000),.out(hidden_layer_out[363:360]));
//Neuron_NN1_layer1 N92 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[44527:44044]),.bias(3'b000),.out(hidden_layer_out[367:364]));
//Neuron_NN1_layer1 N93 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[45011:44528]),.bias(3'b000),.out(hidden_layer_out[371:368]));
//Neuron_NN1_layer1 N94 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[45495:45012]),.bias(3'b000),.out(hidden_layer_out[375:372]));
//Neuron_NN1_layer1 N95 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[45979:45496]),.bias(3'b000),.out(hidden_layer_out[379:376]));
//Neuron_NN1_layer1 N96 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[46463:45980]),.bias(3'b000),.out(hidden_layer_out[383:380]));
//Neuron_NN1_layer1 N97 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[46947:46464]),.bias(3'b000),.out(hidden_layer_out[387:384]));
//Neuron_NN1_layer1 N98 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[47431:46948]),.bias(3'b000),.out(hidden_layer_out[391:388]));
//Neuron_NN1_layer1 N99 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[47915:47432]),.bias(3'b000),.out(hidden_layer_out[395:392]));
//Neuron_NN1_layer1 N100 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[48399:47916]),.bias(3'b000),.out(hidden_layer_out[399:396]));
//Neuron_NN1_layer1 N101 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[48883:48400]),.bias(3'b000),.out(hidden_layer_out[403:400]));
//Neuron_NN1_layer1 N102 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[49367:48884]),.bias(3'b000),.out(hidden_layer_out[407:404]));
//Neuron_NN1_layer1 N103 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[49851:49368]),.bias(3'b000),.out(hidden_layer_out[411:408]));
//Neuron_NN1_layer1 N104 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[50335:49852]),.bias(3'b000),.out(hidden_layer_out[415:412]));
//Neuron_NN1_layer1 N105 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[50819:50336]),.bias(3'b000),.out(hidden_layer_out[419:416]));
//Neuron_NN1_layer1 N106 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[51303:50820]),.bias(3'b000),.out(hidden_layer_out[423:420]));
//Neuron_NN1_layer1 N107 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[51787:51304]),.bias(3'b000),.out(hidden_layer_out[427:424]));
//Neuron_NN1_layer1 N108 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[52271:51788]),.bias(3'b000),.out(hidden_layer_out[431:428]));
//Neuron_NN1_layer1 N109 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[52755:52272]),.bias(3'b000),.out(hidden_layer_out[435:432]));
//Neuron_NN1_layer1 N110 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[53239:52756]),.bias(3'b000),.out(hidden_layer_out[439:436]));
//Neuron_NN1_layer1 N111 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[53723:53240]),.bias(3'b000),.out(hidden_layer_out[443:440]));
//Neuron_NN1_layer1 N112 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[54207:53724]),.bias(3'b000),.out(hidden_layer_out[447:444]));
//Neuron_NN1_layer1 N113 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[54691:54208]),.bias(3'b000),.out(hidden_layer_out[451:448]));
//Neuron_NN1_layer1 N114 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[55175:54692]),.bias(3'b000),.out(hidden_layer_out[455:452]));
//Neuron_NN1_layer1 N115 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[55659:55176]),.bias(3'b000),.out(hidden_layer_out[459:456]));
//Neuron_NN1_layer1 N116 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[56143:55660]),.bias(3'b000),.out(hidden_layer_out[463:460]));
//Neuron_NN1_layer1 N117 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[56627:56144]),.bias(3'b000),.out(hidden_layer_out[467:464]));
//Neuron_NN1_layer1 N118 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[57111:56628]),.bias(3'b000),.out(hidden_layer_out[471:468]));
//Neuron_NN1_layer1 N119 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[57595:57112]),.bias(3'b000),.out(hidden_layer_out[475:472]));
//Neuron_NN1_layer1 N120 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[58079:57596]),.bias(3'b000),.out(hidden_layer_out[479:476]));
//Neuron_NN1_layer1 N121 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[58563:58080]),.bias(3'b000),.out(hidden_layer_out[483:480]));
//Neuron_NN1_layer1 N122 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[59047:58564]),.bias(3'b000),.out(hidden_layer_out[487:484]));
//Neuron_NN1_layer1 N123 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[59531:59048]),.bias(3'b000),.out(hidden_layer_out[491:488]));
//Neuron_NN1_layer1 N124 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[60015:59532]),.bias(3'b000),.out(hidden_layer_out[495:492]));
//Neuron_NN1_layer1 N125 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[60499:60016]),.bias(3'b000),.out(hidden_layer_out[499:496]));
//Neuron_NN1_layer1 N126 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[60983:60500]),.bias(3'b000),.out(hidden_layer_out[503:500]));
//Neuron_NN1_layer1 N127 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[61467:60984]),.bias(3'b000),.out(hidden_layer_out[507:504]));
//Neuron_NN1_layer1 N128 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[61951:61468]),.bias(3'b000),.out(hidden_layer_out[511:508]));
//Neuron_NN1_layer1 N129 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[62435:61952]),.bias(3'b000),.out(hidden_layer_out[515:512]));
//Neuron_NN1_layer1 N130 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[62919:62436]),.bias(3'b000),.out(hidden_layer_out[519:516]));
//Neuron_NN1_layer1 N131 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[63403:62920]),.bias(3'b000),.out(hidden_layer_out[523:520]));
//Neuron_NN1_layer1 N132 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[63887:63404]),.bias(3'b000),.out(hidden_layer_out[527:524]));
//Neuron_NN1_layer1 N133 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[64371:63888]),.bias(3'b000),.out(hidden_layer_out[531:528]));
//Neuron_NN1_layer1 N134 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[64855:64372]),.bias(3'b000),.out(hidden_layer_out[535:532]));
//Neuron_NN1_layer1 N135 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[65339:64856]),.bias(3'b000),.out(hidden_layer_out[539:536]));
//Neuron_NN1_layer1 N136 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[65823:65340]),.bias(3'b000),.out(hidden_layer_out[543:540]));
//Neuron_NN1_layer1 N137 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[66307:65824]),.bias(3'b000),.out(hidden_layer_out[547:544]));
//Neuron_NN1_layer1 N138 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[66791:66308]),.bias(3'b000),.out(hidden_layer_out[551:548]));
//Neuron_NN1_layer1 N139 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[67275:66792]),.bias(3'b000),.out(hidden_layer_out[555:552]));
//Neuron_NN1_layer1 N140 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[67759:67276]),.bias(3'b000),.out(hidden_layer_out[559:556]));
//Neuron_NN1_layer1 N141 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[68243:67760]),.bias(3'b000),.out(hidden_layer_out[563:560]));
//Neuron_NN1_layer1 N142 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[68727:68244]),.bias(3'b000),.out(hidden_layer_out[567:564]));
//Neuron_NN1_layer1 N143 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[69211:68728]),.bias(3'b000),.out(hidden_layer_out[571:568]));
//Neuron_NN1_layer1 N144 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[69695:69212]),.bias(3'b000),.out(hidden_layer_out[575:572]));
//Neuron_NN1_layer1 N145 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[70179:69696]),.bias(3'b000),.out(hidden_layer_out[579:576]));
//Neuron_NN1_layer1 N146 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[70663:70180]),.bias(3'b000),.out(hidden_layer_out[583:580]));
//Neuron_NN1_layer1 N147 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[71147:70664]),.bias(3'b000),.out(hidden_layer_out[587:584]));
//Neuron_NN1_layer1 N148 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[71631:71148]),.bias(3'b000),.out(hidden_layer_out[591:588]));
//Neuron_NN1_layer1 N149 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[72115:71632]),.bias(3'b000),.out(hidden_layer_out[595:592]));
//Neuron_NN1_layer1 N150 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[72599:72116]),.bias(3'b000),.out(hidden_layer_out[599:596]));
//Neuron_NN1_layer1 N151 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[73083:72600]),.bias(3'b000),.out(hidden_layer_out[603:600]));
//Neuron_NN1_layer1 N152 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[73567:73084]),.bias(3'b000),.out(hidden_layer_out[607:604]));
//Neuron_NN1_layer1 N153 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[74051:73568]),.bias(3'b000),.out(hidden_layer_out[611:608]));
//Neuron_NN1_layer1 N154 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[74535:74052]),.bias(3'b000),.out(hidden_layer_out[615:612]));
//Neuron_NN1_layer1 N155 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[75019:74536]),.bias(3'b000),.out(hidden_layer_out[619:616]));
//Neuron_NN1_layer1 N156 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[75503:75020]),.bias(3'b000),.out(hidden_layer_out[623:620]));
//Neuron_NN1_layer1 N157 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[75987:75504]),.bias(3'b000),.out(hidden_layer_out[627:624]));
//Neuron_NN1_layer1 N158 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[76471:75988]),.bias(3'b000),.out(hidden_layer_out[631:628]));
//Neuron_NN1_layer1 N159 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[76955:76472]),.bias(3'b000),.out(hidden_layer_out[635:632]));
//Neuron_NN1_layer1 N160 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[77439:76956]),.bias(3'b000),.out(hidden_layer_out[639:636]));
//Neuron_NN1_layer1 N161 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[77923:77440]),.bias(3'b000),.out(hidden_layer_out[643:640]));
//Neuron_NN1_layer1 N162 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[78407:77924]),.bias(3'b000),.out(hidden_layer_out[647:644]));
//Neuron_NN1_layer1 N163 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[78891:78408]),.bias(3'b000),.out(hidden_layer_out[651:648]));
//Neuron_NN1_layer1 N164 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[79375:78892]),.bias(3'b000),.out(hidden_layer_out[655:652]));
//Neuron_NN1_layer1 N165 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[79859:79376]),.bias(3'b000),.out(hidden_layer_out[659:656]));
//Neuron_NN1_layer1 N166 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[80343:79860]),.bias(3'b000),.out(hidden_layer_out[663:660]));
//Neuron_NN1_layer1 N167 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[80827:80344]),.bias(3'b000),.out(hidden_layer_out[667:664]));
//Neuron_NN1_layer1 N168 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[81311:80828]),.bias(3'b000),.out(hidden_layer_out[671:668]));
//Neuron_NN1_layer1 N169 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[81795:81312]),.bias(3'b000),.out(hidden_layer_out[675:672]));
//Neuron_NN1_layer1 N170 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[82279:81796]),.bias(3'b000),.out(hidden_layer_out[679:676]));
//Neuron_NN1_layer1 N171 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[82763:82280]),.bias(3'b000),.out(hidden_layer_out[683:680]));
//Neuron_NN1_layer1 N172 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[83247:82764]),.bias(3'b000),.out(hidden_layer_out[687:684]));
//Neuron_NN1_layer1 N173 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[83731:83248]),.bias(3'b000),.out(hidden_layer_out[691:688]));
//Neuron_NN1_layer1 N174 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[84215:83732]),.bias(3'b000),.out(hidden_layer_out[695:692]));
//Neuron_NN1_layer1 N175 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[84699:84216]),.bias(3'b000),.out(hidden_layer_out[699:696]));
//Neuron_NN1_layer1 N176 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[85183:84700]),.bias(3'b000),.out(hidden_layer_out[703:700]));
//Neuron_NN1_layer1 N177 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[85667:85184]),.bias(3'b000),.out(hidden_layer_out[707:704]));
//Neuron_NN1_layer1 N178 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[86151:85668]),.bias(3'b000),.out(hidden_layer_out[711:708]));
//Neuron_NN1_layer1 N179 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[86635:86152]),.bias(3'b000),.out(hidden_layer_out[715:712]));
//Neuron_NN1_layer1 N180 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[87119:86636]),.bias(3'b000),.out(hidden_layer_out[719:716]));
//Neuron_NN1_layer1 N181 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[87603:87120]),.bias(3'b000),.out(hidden_layer_out[723:720]));
//Neuron_NN1_layer1 N182 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[88087:87604]),.bias(3'b000),.out(hidden_layer_out[727:724]));
//Neuron_NN1_layer1 N183 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[88571:88088]),.bias(3'b000),.out(hidden_layer_out[731:728]));
//Neuron_NN1_layer1 N184 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[89055:88572]),.bias(3'b000),.out(hidden_layer_out[735:732]));
//Neuron_NN1_layer1 N185 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[89539:89056]),.bias(3'b000),.out(hidden_layer_out[739:736]));
//Neuron_NN1_layer1 N186 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[90023:89540]),.bias(3'b000),.out(hidden_layer_out[743:740]));
//Neuron_NN1_layer1 N187 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[90507:90024]),.bias(3'b000),.out(hidden_layer_out[747:744]));
//Neuron_NN1_layer1 N188 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[90991:90508]),.bias(3'b000),.out(hidden_layer_out[751:748]));
//Neuron_NN1_layer1 N189 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[91475:90992]),.bias(3'b000),.out(hidden_layer_out[755:752]));
//Neuron_NN1_layer1 N190 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[91959:91476]),.bias(3'b000),.out(hidden_layer_out[759:756]));
//Neuron_NN1_layer1 N191 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[92443:91960]),.bias(3'b000),.out(hidden_layer_out[763:760]));
//Neuron_NN1_layer1 N192 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[92927:92444]),.bias(3'b000),.out(hidden_layer_out[767:764]));
//Neuron_NN1_layer1 N193 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[93411:92928]),.bias(3'b000),.out(hidden_layer_out[771:768]));
//Neuron_NN1_layer1 N194 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[93895:93412]),.bias(3'b000),.out(hidden_layer_out[775:772]));
//Neuron_NN1_layer1 N195 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[94379:93896]),.bias(3'b000),.out(hidden_layer_out[779:776]));
//Neuron_NN1_layer1 N196 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[94863:94380]),.bias(3'b000),.out(hidden_layer_out[783:780]));
//Neuron_NN1_layer1 N197 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[95347:94864]),.bias(3'b000),.out(hidden_layer_out[787:784]));
//Neuron_NN1_layer1 N198 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[95831:95348]),.bias(3'b000),.out(hidden_layer_out[791:788]));
//Neuron_NN1_layer1 N199 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[96315:95832]),.bias(3'b000),.out(hidden_layer_out[795:792]));
//Neuron_NN1_layer1 N200 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[96799:96316]),.bias(3'b000),.out(hidden_layer_out[799:796]));

Neuron_NN1_layer1 N1 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[483:0]),.bias(3'b000),.out(hidden_layer_out[3:0]));
Neuron_NN1_layer1 N2 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[967:484]),.bias(3'b000),.out(hidden_layer_out[7:4]));
Neuron_NN1_layer1 N3 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[1451:968]),.bias(3'b000),.out(hidden_layer_out[11:8]));
Neuron_NN1_layer1 N4 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[1935:1452]),.bias(3'b000),.out(hidden_layer_out[15:12]));
Neuron_NN1_layer1 N5 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[2419:1936]),.bias(3'b000),.out(hidden_layer_out[19:16]));
Neuron_NN1_layer1 N6 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[2903:2420]),.bias(3'b000),.out(hidden_layer_out[23:20]));
Neuron_NN1_layer1 N7 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[3387:2904]),.bias(3'b000),.out(hidden_layer_out[27:24]));
Neuron_NN1_layer1 N8 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[3871:3388]),.bias(3'b000),.out(hidden_layer_out[31:28]));
Neuron_NN1_layer1 N9 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[4355:3872]),.bias(3'b000),.out(hidden_layer_out[35:32]));
Neuron_NN1_layer1 N10 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[4839:4356]),.bias(3'b000),.out(hidden_layer_out[39:36]));
Neuron_NN1_layer1 N11 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[5323:4840]),.bias(3'b000),.out(hidden_layer_out[43:40]));
Neuron_NN1_layer1 N12 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[5807:5324]),.bias(3'b000),.out(hidden_layer_out[47:44]));
Neuron_NN1_layer1 N13 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[6291:5808]),.bias(3'b000),.out(hidden_layer_out[51:48]));
Neuron_NN1_layer1 N14 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[6775:6292]),.bias(3'b000),.out(hidden_layer_out[55:52]));
Neuron_NN1_layer1 N15 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[7259:6776]),.bias(3'b000),.out(hidden_layer_out[59:56]));
Neuron_NN1_layer1 N16 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[7743:7260]),.bias(3'b000),.out(hidden_layer_out[63:60]));
Neuron_NN1_layer1 N17 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[8227:7744]),.bias(3'b000),.out(hidden_layer_out[67:64]));
Neuron_NN1_layer1 N18 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[8711:8228]),.bias(3'b000),.out(hidden_layer_out[71:68]));
Neuron_NN1_layer1 N19 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[9195:8712]),.bias(3'b000),.out(hidden_layer_out[75:72]));
Neuron_NN1_layer1 N20 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[9679:9196]),.bias(3'b000),.out(hidden_layer_out[79:76]));
Neuron_NN1_layer1 N21 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[10163:9680]),.bias(3'b000),.out(hidden_layer_out[83:80]));
Neuron_NN1_layer1 N22 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[10647:10164]),.bias(3'b000),.out(hidden_layer_out[87:84]));
Neuron_NN1_layer1 N23 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[11131:10648]),.bias(3'b000),.out(hidden_layer_out[91:88]));
Neuron_NN1_layer1 N24 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[11615:11132]),.bias(3'b000),.out(hidden_layer_out[95:92]));
Neuron_NN1_layer1 N25 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[12099:11616]),.bias(3'b000),.out(hidden_layer_out[99:96]));
Neuron_NN1_layer1 N26 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[12583:12100]),.bias(3'b000),.out(hidden_layer_out[103:100]));
Neuron_NN1_layer1 N27 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[13067:12584]),.bias(3'b000),.out(hidden_layer_out[107:104]));
Neuron_NN1_layer1 N28 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[13551:13068]),.bias(3'b000),.out(hidden_layer_out[111:108]));
Neuron_NN1_layer1 N29 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[14035:13552]),.bias(3'b000),.out(hidden_layer_out[115:112]));
Neuron_NN1_layer1 N30 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[14519:14036]),.bias(3'b000),.out(hidden_layer_out[119:116]));
Neuron_NN1_layer1 N31 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[15003:14520]),.bias(3'b000),.out(hidden_layer_out[123:120]));
Neuron_NN1_layer1 N32 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[15487:15004]),.bias(3'b000),.out(hidden_layer_out[127:124]));
Neuron_NN1_layer1 N33 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[15971:15488]),.bias(3'b000),.out(hidden_layer_out[131:128]));
Neuron_NN1_layer1 N34 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[16455:15972]),.bias(3'b000),.out(hidden_layer_out[135:132]));
Neuron_NN1_layer1 N35 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[16939:16456]),.bias(3'b000),.out(hidden_layer_out[139:136]));
Neuron_NN1_layer1 N36 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[17423:16940]),.bias(3'b000),.out(hidden_layer_out[143:140]));
Neuron_NN1_layer1 N37 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[17907:17424]),.bias(3'b000),.out(hidden_layer_out[147:144]));
Neuron_NN1_layer1 N38 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[18391:17908]),.bias(3'b000),.out(hidden_layer_out[151:148]));
Neuron_NN1_layer1 N39 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[18875:18392]),.bias(3'b000),.out(hidden_layer_out[155:152]));
Neuron_NN1_layer1 N40 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[19359:18876]),.bias(3'b000),.out(hidden_layer_out[159:156]));
Neuron_NN1_layer1 N41 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[19843:19360]),.bias(3'b000),.out(hidden_layer_out[163:160]));
Neuron_NN1_layer1 N42 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[20327:19844]),.bias(3'b000),.out(hidden_layer_out[167:164]));
Neuron_NN1_layer1 N43 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[20811:20328]),.bias(3'b000),.out(hidden_layer_out[171:168]));
Neuron_NN1_layer1 N44 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[21295:20812]),.bias(3'b000),.out(hidden_layer_out[175:172]));
Neuron_NN1_layer1 N45 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[21779:21296]),.bias(3'b000),.out(hidden_layer_out[179:176]));
Neuron_NN1_layer1 N46 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[22263:21780]),.bias(3'b000),.out(hidden_layer_out[183:180]));
Neuron_NN1_layer1 N47 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[22747:22264]),.bias(3'b000),.out(hidden_layer_out[187:184]));
Neuron_NN1_layer1 N48 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[23231:22748]),.bias(3'b000),.out(hidden_layer_out[191:188]));
Neuron_NN1_layer1 N49 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[23715:23232]),.bias(3'b000),.out(hidden_layer_out[195:192]));
Neuron_NN1_layer1 N50 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[24199:23716]),.bias(3'b000),.out(hidden_layer_out[199:196]));
Neuron_NN1_layer1 N51 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[24683:24200]),.bias(3'b000),.out(hidden_layer_out[203:200]));
Neuron_NN1_layer1 N52 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[25167:24684]),.bias(3'b000),.out(hidden_layer_out[207:204]));
Neuron_NN1_layer1 N53 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[25651:25168]),.bias(3'b000),.out(hidden_layer_out[211:208]));
Neuron_NN1_layer1 N54 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[26135:25652]),.bias(3'b000),.out(hidden_layer_out[215:212]));
Neuron_NN1_layer1 N55 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[26619:26136]),.bias(3'b000),.out(hidden_layer_out[219:216]));
Neuron_NN1_layer1 N56 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[27103:26620]),.bias(3'b000),.out(hidden_layer_out[223:220]));
Neuron_NN1_layer1 N57 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[27587:27104]),.bias(3'b000),.out(hidden_layer_out[227:224]));
Neuron_NN1_layer1 N58 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[28071:27588]),.bias(3'b000),.out(hidden_layer_out[231:228]));
Neuron_NN1_layer1 N59 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[28555:28072]),.bias(3'b000),.out(hidden_layer_out[235:232]));
Neuron_NN1_layer1 N60 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[29039:28556]),.bias(3'b000),.out(hidden_layer_out[239:236]));
Neuron_NN1_layer1 N61 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[29523:29040]),.bias(3'b000),.out(hidden_layer_out[243:240]));
Neuron_NN1_layer1 N62 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[30007:29524]),.bias(3'b000),.out(hidden_layer_out[247:244]));
Neuron_NN1_layer1 N63 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[30491:30008]),.bias(3'b000),.out(hidden_layer_out[251:248]));
Neuron_NN1_layer1 N64 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[30975:30492]),.bias(3'b000),.out(hidden_layer_out[255:252]));
Neuron_NN1_layer1 N65 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[31459:30976]),.bias(3'b000),.out(hidden_layer_out[259:256]));
Neuron_NN1_layer1 N66 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[31943:31460]),.bias(3'b000),.out(hidden_layer_out[263:260]));
Neuron_NN1_layer1 N67 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[32427:31944]),.bias(3'b000),.out(hidden_layer_out[267:264]));
Neuron_NN1_layer1 N68 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[32911:32428]),.bias(3'b000),.out(hidden_layer_out[271:268]));
Neuron_NN1_layer1 N69 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[33395:32912]),.bias(3'b000),.out(hidden_layer_out[275:272]));
Neuron_NN1_layer1 N70 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[33879:33396]),.bias(3'b000),.out(hidden_layer_out[279:276]));
Neuron_NN1_layer1 N71 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[34363:33880]),.bias(3'b000),.out(hidden_layer_out[283:280]));
Neuron_NN1_layer1 N72 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[34847:34364]),.bias(3'b000),.out(hidden_layer_out[287:284]));
Neuron_NN1_layer1 N73 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[35331:34848]),.bias(3'b000),.out(hidden_layer_out[291:288]));
Neuron_NN1_layer1 N74 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[35815:35332]),.bias(3'b000),.out(hidden_layer_out[295:292]));
Neuron_NN1_layer1 N75 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[36299:35816]),.bias(3'b000),.out(hidden_layer_out[299:296]));
Neuron_NN1_layer1 N76 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[36783:36300]),.bias(3'b000),.out(hidden_layer_out[303:300]));
Neuron_NN1_layer1 N77 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[37267:36784]),.bias(3'b000),.out(hidden_layer_out[307:304]));
Neuron_NN1_layer1 N78 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[37751:37268]),.bias(3'b000),.out(hidden_layer_out[311:308]));
Neuron_NN1_layer1 N79 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[38235:37752]),.bias(3'b000),.out(hidden_layer_out[315:312]));
Neuron_NN1_layer1 N80 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[38719:38236]),.bias(3'b000),.out(hidden_layer_out[319:316]));
Neuron_NN1_layer1 N81 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[39203:38720]),.bias(3'b000),.out(hidden_layer_out[323:320]));
Neuron_NN1_layer1 N82 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[39687:39204]),.bias(3'b000),.out(hidden_layer_out[327:324]));
Neuron_NN1_layer1 N83 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[40171:39688]),.bias(3'b000),.out(hidden_layer_out[331:328]));
Neuron_NN1_layer1 N84 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[40655:40172]),.bias(3'b000),.out(hidden_layer_out[335:332]));
Neuron_NN1_layer1 N85 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[41139:40656]),.bias(3'b000),.out(hidden_layer_out[339:336]));
Neuron_NN1_layer1 N86 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[41623:41140]),.bias(3'b000),.out(hidden_layer_out[343:340]));
Neuron_NN1_layer1 N87 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[42107:41624]),.bias(3'b000),.out(hidden_layer_out[347:344]));
Neuron_NN1_layer1 N88 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[42591:42108]),.bias(3'b000),.out(hidden_layer_out[351:348]));
Neuron_NN1_layer1 N89 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[43075:42592]),.bias(3'b000),.out(hidden_layer_out[355:352]));
Neuron_NN1_layer1 N90 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[43559:43076]),.bias(3'b000),.out(hidden_layer_out[359:356]));
Neuron_NN1_layer1 N91 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[44043:43560]),.bias(3'b000),.out(hidden_layer_out[363:360]));
Neuron_NN1_layer1 N92 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[44527:44044]),.bias(3'b000),.out(hidden_layer_out[367:364]));
Neuron_NN1_layer1 N93 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[45011:44528]),.bias(3'b000),.out(hidden_layer_out[371:368]));
Neuron_NN1_layer1 N94 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[45495:45012]),.bias(3'b000),.out(hidden_layer_out[375:372]));
Neuron_NN1_layer1 N95 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[45979:45496]),.bias(3'b000),.out(hidden_layer_out[379:376]));
Neuron_NN1_layer1 N96 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[46463:45980]),.bias(3'b000),.out(hidden_layer_out[383:380]));
Neuron_NN1_layer1 N97 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[46947:46464]),.bias(3'b000),.out(hidden_layer_out[387:384]));
Neuron_NN1_layer1 N98 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[47431:46948]),.bias(3'b000),.out(hidden_layer_out[391:388]));
Neuron_NN1_layer1 N99 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[47915:47432]),.bias(3'b000),.out(hidden_layer_out[395:392]));
Neuron_NN1_layer1 N100 (.reset2(reset2),.clk3(clk3),.input_features(input_features),.input_weights(weights_NN1_layer1[48399:47916]),.bias(3'b000),.out(hidden_layer_out[399:396]));

 
//////////////////////////////Output Layer 10 Nodes/////////////////////////////////////// 

// NN1(.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[119:0]),.bias(3'b000),.out(output_layer_out[0])); 
//Neuron_NN1_layer2 NN2 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[239:120]),.bias(3'b000),.out(output_layer_out[1]));
//Neuron_NN1_layer2 NN3 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[359:240]),.bias(3'b000),.out(output_layer_out[2]));
//Neuron_NN1_layer2 NN4 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[479:360]),.bias(3'b000),.out(output_layer_out[3]));
//Neuron_NN1_layer2 NN5 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[599:480]),.bias(3'b000),.out(output_layer_out[4]));
//Neuron_NN1_layer2 NN6 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[719:600]),.bias(3'b000),.out(output_layer_out[5]));
//Neuron_NN1_layer2 NN7 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[839:720]),.bias(3'b000),.out(output_layer_out[6]));
//Neuron_NN1_layer2 NN8 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[959:840]),.bias(3'b000),.out(output_layer_out[7]));
//Neuron_NN1_layer2 NN9 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[1079:960]),.bias(3'b000),.out(output_layer_out[8]));
//Neuron_NN1_layer2 NN10 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[1199:1080]),.bias(3'b000),.out(output_layer_out[9]));

Neuron_NN1_layer2 NN1(.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[399:0]),.bias(3'b000),.out(output_layer_out[0])); 
Neuron_NN1_layer2 NN2 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[799:400]),.bias(3'b000),.out(output_layer_out[1]));
Neuron_NN1_layer2 NN3 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[1199:800]),.bias(3'b000),.out(output_layer_out[2]));
Neuron_NN1_layer2 NN4 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[1599:1200]),.bias(3'b000),.out(output_layer_out[3]));
Neuron_NN1_layer2 NN5 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[1999:1600]),.bias(3'b000),.out(output_layer_out[4]));
Neuron_NN1_layer2 NN6 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[2399:2000]),.bias(3'b000),.out(output_layer_out[5]));
Neuron_NN1_layer2 NN7 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[2799:2400]),.bias(3'b000),.out(output_layer_out[6]));
Neuron_NN1_layer2 NN8 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[3199:2800]),.bias(3'b000),.out(output_layer_out[7]));
Neuron_NN1_layer2 NN9 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[3599:3200]),.bias(3'b000),.out(output_layer_out[8]));
Neuron_NN1_layer2 NN10 (.reset1(reset2),.clk3(clk3),.input_features(hidden_layer_out),.input_weights(weights_NN1_layer2[3999:3600]),.bias(3'b000),.out(output_layer_out[9]));




/////////////////////////////Get the final output by looking at the highest value for "output_layer_out"/////////////////////////////////////////////////////////




always @(output_layer_out[0] or output_layer_out[1] or output_layer_out[2] or output_layer_out[3] or output_layer_out[4] or output_layer_out[5] or output_layer_out[6] or output_layer_out[7] or output_layer_out[8] or output_layer_out[9])
begin

if (output_layer_out[0] >= output_layer_out[1])begin
max=output_layer_out[0];
final_output=0;end
else begin
max=output_layer_out[1];
final_output=1;end

if (output_layer_out[2]>max) begin
max=output_layer_out[2];
final_output=2;end

if (output_layer_out[3]>max)begin
max=output_layer_out[3];
final_output=3;end

if (output_layer_out[4]>max)begin
max=output_layer_out[4];
final_output=4;end

if (output_layer_out[5]>max)begin
max=output_layer_out[5];
final_output=5;end

if (output_layer_out[6]>max)begin
max=output_layer_out[6];
final_output=6;end

if (output_layer_out[7]>max)begin
max=output_layer_out[7];
final_output=7;end

if (output_layer_out[8]>max)begin
max=output_layer_out[8];
final_output=8;end

if (output_layer_out[9]>max)begin
max=output_layer_out[9];
final_output=9;end

end


input_rx U2(
.clk(clk)     , // Top level system clock input.
.sw_0(sw_0)    , // Slide switches.
.rst(rst),
//input               sw_1    , // Slide switches.
.uart_rxd(uart_rxd), // UART Recieve pin.
.input_valid(led1),
//output  wire        uart_txd, // UART transmit pin.
//output wire [127:0] led2,
.network_input(input_features0)
);

clk_div_n #(
.WIDTH(WIDTH)) i_clk_div_n(
.clk(clk),
.reset(1'b0),
.div_num(div_num),
.clk_out(clk3)
);

// signals
    wire [9:0] w_x, w_y;
    wire w_video_on, w_p_tick;
    reg [11:0] rgb_reg;
    wire [11:0] rgb_next;


    // VGA Controller
    vga_controller vga(.clk_100MHz(clk), .reset(reset), .hsync(hsync), .vsync(vsync),
                       .video_on(w_video_on), .p_tick(w_p_tick), .x(w_x), .y(w_y));
//    // Text Generation Circuit
    ascii_test at(.clk(clk), .video_on(w_video_on), .x(w_x), .y(w_y), .rgb(rgb_next), .reset2(reset2), .SW(final_output1), .a_to_g(a_to_g), .rst(rst), .an(AN), .dp(DP), .BTNR(BTNR));

//    // rgb buffer
    always @(posedge clk)
        if(w_p_tick)
            rgb_reg <= rgb_next;
            
//    // output
    assign rgb = rgb_reg;
endmodule